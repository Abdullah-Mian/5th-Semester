library ieee;
use ieee.std_logic_1164.all;

package MyPackage is
    component Dflipflop is
        port (
            clk   : in std_logic;
            D     : in std_logic;
            Q     : out std_logic;
            Qnot  : out std_logic
        );
    end component;
end package MyPackage;